`timescale 1ns / 1ps

module cla32
(
    input wire[31:0] a,
    input wire[31:0] b,
    input wire cin,
    output wire cout,
    output wire[31:0] sum
);

genvar i;
wire[31:0] carry;

// Carry Generation
assign carry[0]  = cin;
assign carry[1]  = (a[0] & b[0])   | ((a[0] ^ b[0])   & cin);
assign carry[2]  = (a[1] & b[1])   | ((a[1] ^ b[1])   & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))));
assign carry[3]  = (a[2] & b[2])   | ((a[2] ^ b[2])   & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))));
assign carry[4]  = (a[3] & b[3])   | ((a[3] ^ b[3])   & ((a[2] & b[2])   | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))));
assign carry[5]  = (a[4] & b[4])   | ((a[4] ^ b[4])   & ((a[3] & b[3])   | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))));
assign carry[6]  = (a[5] & b[5])   | ((a[5] ^ b[5])   & ((a[4] & b[4])   | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))));
assign carry[7]  = (a[6] & b[6])   | ((a[6] ^ b[6])   & ((a[5] & b[5])   | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))));
assign carry[8]  = (a[7] & b[7])   | ((a[7] ^ b[7])   & ((a[6] & b[6])   | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))));
assign carry[9]  = (a[8] & b[8])   | ((a[8] ^ b[8])   & ((a[7] & b[7])   | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))));
assign carry[10] = (a[9] & b[9])   | ((a[9] ^ b[9])   & ((a[8] & b[8])   | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))));
assign carry[11] = (a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))));
assign carry[12] = (a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))));
assign carry[13] = (a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))));
assign carry[14] = (a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))));
assign carry[15] = (a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))));
assign carry[16] = (a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))));
assign carry[17] = (a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))));
assign carry[18] = (a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))));
assign carry[19] = (a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))));
assign carry[20] = (a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))));
assign carry[21] = (a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))));
assign carry[22] = (a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))));
assign carry[23] = (a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])    | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))));
assign carry[24] = (a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])     | ((a[1] ^ b[1]) & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))));
assign carry[25] = (a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])     | ((a[2] ^ b[2]) & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))))));
assign carry[26] = (a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])     | ((a[3] ^ b[3]) & ((a[2] & b[2])   | ((a[2] ^ b[2]) & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))))))));
assign carry[27] = (a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])     | ((a[4] ^ b[4]) & ((a[3] & b[3])   | ((a[3] ^ b[3]) & ((a[2] & b[2])   | ((a[2] ^ b[2]) & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))))))))));
assign carry[28] = (a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])     | ((a[5] ^ b[5]) & ((a[4] & b[4])   | ((a[4] ^ b[4]) & ((a[3] & b[3])   | ((a[3] ^ b[3]) & ((a[2] & b[2])   | ((a[2] ^ b[2]) & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))))))))))));
assign carry[29] = (a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])     | ((a[6] ^ b[6]) & ((a[5] & b[5])   | ((a[5] ^ b[5]) & ((a[4] & b[4])   | ((a[4] ^ b[4]) & ((a[3] & b[3])   | ((a[3] ^ b[3]) & ((a[2] & b[2])   | ((a[2] ^ b[2]) & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
assign carry[30] = (a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])     | ((a[7] ^ b[7]) & ((a[6] & b[6])   | ((a[6] ^ b[6]) & ((a[5] & b[5])   | ((a[5] ^ b[5]) & ((a[4] & b[4])   | ((a[4] ^ b[4]) & ((a[3] & b[3])   | ((a[3] ^ b[3]) & ((a[2] & b[2])   | ((a[2] ^ b[2]) & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
assign carry[31] = (a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])     | ((a[8] ^ b[8]) & ((a[7] & b[7])   | ((a[7] ^ b[7]) & ((a[6] & b[6])   | ((a[6] ^ b[6]) & ((a[5] & b[5])   | ((a[5] ^ b[5]) & ((a[4] & b[4])   | ((a[4] ^ b[4]) & ((a[3] & b[3])   | ((a[3] ^ b[3]) & ((a[2] & b[2])   | ((a[2] ^ b[2]) & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0])  | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
assign cout      = (a[31] & b[31]) | ((a[31] ^ b[31]) & ((a[30] & b[30]) | ((a[30] ^ b[30]) & ((a[29] & b[29]) | ((a[29] ^ b[29]) & ((a[28] & b[28]) | ((a[28] ^ b[28]) & ((a[27] & b[27]) | ((a[27] ^ b[27]) & ((a[26] & b[26]) | ((a[26] ^ b[26]) & ((a[25] & b[25]) | ((a[25] ^ b[25]) & ((a[24] & b[24]) | ((a[24] ^ b[24]) & ((a[23] & b[23]) | ((a[23] ^ b[23]) & ((a[22] & b[22]) | ((a[22] ^ b[22]) & ((a[21] & b[21]) | ((a[21] ^ b[21]) & ((a[20] & b[20]) | ((a[20] ^ b[20]) & ((a[19] & b[19]) | ((a[19] ^ b[19]) & ((a[18] & b[18]) | ((a[18] ^ b[18]) & ((a[17] & b[17]) | ((a[17] ^ b[17]) & ((a[16] & b[16]) | ((a[16] ^ b[16]) & ((a[15] & b[15]) | ((a[15] ^ b[15]) & ((a[14] & b[14]) | ((a[14] ^ b[14]) & ((a[13] & b[13]) | ((a[13] ^ b[13]) & ((a[12] & b[12]) | ((a[12] ^ b[12]) & ((a[11] & b[11]) | ((a[11] ^ b[11]) & ((a[10] & b[10]) | ((a[10] ^ b[10]) & ((a[9] & b[9])   | ((a[9] ^ b[9]) & ((a[8] & b[8])   | ((a[8] ^ b[8]) & ((a[7] & b[7])   | ((a[7] ^ b[7]) & ((a[6] & b[6])   | ((a[6] ^ b[6]) & ((a[5] & b[5])   | ((a[5] ^ b[5]) & ((a[4] & b[4])   | ((a[4] ^ b[4]) & ((a[3] & b[3])   | ((a[3] ^ b[3]) & ((a[2] & b[2])   | ((a[2] ^ b[2]) & ((a[1] & b[1])   | ((a[1] ^ b[1]) & (((a[0] & b[0]) | ((a[0] ^ b[0]) & cin))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));


// Generate Adders
generate
    for (i = 0; i < 32; i = i + 1)
    begin
        full_adder gen_add
        (
            .a(a[i]),
            .b(b[i]),
            .cin(carry[i]),
            .s(sum[i]),
            .cout()
        );
    end
endgenerate

endmodule
